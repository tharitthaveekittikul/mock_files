This is a mock file for file_621.vhd