This is a mock file for file_306.vhd