This is a mock file for file_486.vhd