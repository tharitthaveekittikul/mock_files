This is a mock file for file_512.vhd