This is a mock file for file_497.vhd