This is a mock file for file_179.vhd