This is a mock file for file_550.vhd